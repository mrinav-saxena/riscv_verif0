class cache_env ;



endclass : cache_env

class cache_test ;

    cache_env env_inst ;
    cache_if cache_if_inst ;


endclass : cache_test