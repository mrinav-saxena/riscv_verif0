interface cache_if () ;

endinterface : cache_if